LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.all;

ENTITY DDS IS
PORT(CLOCK_50:IN STD_LOGIC;
	  KEY: IN STD_LOGIC_VECTOR(3 DOWNTO 0);	    --input to change the frequency sweep
     GPIO: INOUT STD_LOGIC_VECTOR (8 DOWNTO 0));    --Output to the DAC
END DDS;

ARCHITECTURE RTL OF DDS IS

COMPONENT ROM IS                                        --Port map to the ROM
PORT (
		address	 : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		clock: IN STD_LOGIC;
		q: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END COMPONENT;
SIGNAL ACC:INTEGER:=0;
SIGNAL PI:INTEGER :=1000;

SIGNAL TEMP:STD_LOGIC_VECTOR (31 DOWNTO 0);
SIGNAL ADDRESS:STD_LOGIC_VECTOR (5 DOWNTO 0);
SIGNAL DATA_T: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL COUNTER : STD_LOGIC_VECTOR(12 DOWNTO 0);
SIGNAL TEMP_DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL TICK: INTEGER RANGE 0 TO 11:= 1;
SIGNAL COUNT: INTEGER RANGE 1 TO 20833:=1;
SIGNAL TRIGGER: STD_LOGIC;
SIGNAL DPI: INTEGER:=2828;
SIGNAL DFDT: INTEGER:= 4;
SIGNAL DFDT0,DFDT1,DFDT2,DFDT3:INTEGER:=0;
SIGNAL DATAOUT:STD_LOGIC_VECTOR(7 DOWNTO 0);
CONSTANT CONST: REAL:= 0.282;
SIGNAL STATE:STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN

rom_inst : rom PORT MAP (address	 => ADDRESS,clock	 => CLOCK_50,q	 => TEMP_DATA);
PROCESS(TEMP_DATA)                                             --Handles the convertion of 8 bit to 6 bit look up table
BEGIN
	CASE STATE IS
		WHEN "00"=> DATAOUT<=std_logic_vector(to_unsigned(to_integer(unsigned(TEMP_DATA)),8));
		WHEN "01"=> DATAOUT<=std_logic_vector(to_unsigned(to_integer(unsigned(TEMP_DATA)),8));
		WHEN "10"=> DATAOUT<=std_logic_vector(to_unsigned(255-to_integer(unsigned(TEMP_DATA)),8));
		WHEN "11"=> DATAOUT<=std_logic_vector(to_unsigned(255-to_integer(unsigned(TEMP_DATA)),8));
	END CASE;
END PROCESS;
GPIO(7 downto 0)<=DATAOUT;
PROCESS(TEMP)
BEGIN
	IF (TEMP>="00000000" AND TEMP<"01000000") THEN
		ADDRESS<=TEMP(5 DOWNTO 0);
		STATE<="00";
	ELSIF (TEMP>="01000000" AND TEMP<"10000000") THEN
		ADDRESS<=(not TEMP(5 DOWNTO 0));
		STATE<="01";
	ELSIF (TEMP>="10000000" AND TEMP<"11000000") THEN
		ADDRESS<=TEMP(5 DOWNTO 0);
		STATE<="10";
	ELSE 
		ADDRESS<=(not TEMP(5 DOWNTO 0));
		STATE<="11";
	END IF;
END PROCESS;

PROCESS(CLOCK_50)             --clock divider for the Sampling rate
BEGIN
IF(rising_edge(CLOCK_50)) THEN
TICK<=TICK+1;
IF(TICK=2) THEN
GPIO(8)<=GPIO(8) XOR '1';
TICK<=1;
END IF;
END IF;
END PROCESS;

PROCESS(TICK,GPIO(8))             
BEGIN
IF (rising_edge(GPIO(8))) THEN
ACC<=ACC+PI;
TEMP<=STD_LOGIC_VECTOR(TO_UNSIGNED(ACC,32));
END IF;
END PROCESS;

PROCESS(CLOCK_50)              --clock divider for the changing PI
BEGIN
IF(rising_edge(CLOCK_50)) THEN
COUNT<=COUNT+1;
IF(COUNT = 20833) THEN
TRIGGER <= TRIGGER XOR '1';
COUNT <= 1;
END IF;
END IF;
END PROCESS;

PROCESS(TRIGGER)      --actual adding of PI to change frequency
BEGIN
IF(rising_edge(TRIGGER)) THEN
PI <= PI + DPI;
IF(PI > 138006897 ) THEN
PI <= 1;
END IF;
END IF;
END PROCESS;

PROCESS(KEY)
BEGIN

IF(RISing_edge(KEY(0))) THEN
DFDT0 <= DFDT0 + 1;
END IF;
IF(RISing_edge(KEY(1))) THEN
DFDT1 <= DFDT1 + 10;
END IF;
IF(RISing_edge(KEY(2))) THEN
DFDT2 <= DFDT2 + 100;
END IF;
IF(RISing_edge(KEY(3))) THEN
DFDT3 <= DFDT3 + 1000;
END IF;
DFDT<=DFDT0+DFDT1+DFDT2+DFDT3;
DPI<=INTEGER(282*DFDT/1000);
IF(DFDT > 14500) THEN
DFDT <= 14500;
END IF;
END PROCESS;


END RTL;	
